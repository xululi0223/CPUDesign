module decoder_5_32(
    input  [ 4:0] in,
    output [31:0] out
);

genvar i;
generate for (i=0; i<32; i=i+1) begin : gen_for_dec_5_32
    assign out[i] = (in == i);
end endgenerate

endmodule


module decoder_6_64(
    input  [ 5:0] in,
    output [63:0] out
);

genvar i;
/**************修改***************/
generate for (i=0; i<64; i=i+1) begin : gen_for_dec_6_64 //generate for (i=0; i<63; i=i+1) begin : gen_for_dec_6_64 源代码 应该是i<64
/**************修改完毕***************/
    assign out[i] = (in == i);
end endgenerate

endmodule

